`timescale 1ns / 1ps

/* �����֮�ǡ� */
module song3(clk_5MHz,clk_4Hz,select,beep);
	
input clk_5MHz,clk_4Hz,select;			
output beep;					  

reg  [3:0]high,med,low;
reg  [15:0]origin;
reg	beep_r;					  
reg  [7:0]state;					
reg  [15:0]count;			

assign beep = beep_r;	     

/* �������������� */
always @(posedge clk_5MHz)
begin
	/* ������ */
	count <= count + 1'b1;		
	if(count == origin)
	begin
		/* ���������� */
		count <= 16'h0;			
		/* ���ȡ�� */
		beep_r <= !beep_r;		
	end
end

/* �������ת�� */
always@(posedge clk_4Hz)
begin
	if(select)
	begin
		case({high,med,low})
			'b000000000001:origin=22900; //��1
			'b000000000010:origin=20408; //��2
			'b000000000011:origin=18181; //��3
			'b000000000100:origin=17142; //��4
			'b000000000101:origin=15267; //��5
			'b000000000110:origin=13605; //��6
			'b000000000111:origin=12121; //��7
			'b000000010000:origin=11472; //��1
			'b000000100000:origin=10216; //��2
			'b000000110000:origin=9101;  //��3
			'b000000111000:origin=8571;  //��4
			'b000001010000:origin=7653;  //��5
			'b000001100000:origin=6818;  //��6
			'b000010000000:origin=6060;  //��7
			'b000100000000:origin=5733;  //��1
			'b001000000000:origin=5108;  //��2
			'b001100000000:origin=4551;  //��3
			'b001010000000:origin=4294;  //��4
			'b010000000000:origin=3826;  //��5
			'b011000000000:origin=3409;  //��6
			'b010100000000:origin=3050;  //��7
		endcase
	end
	
	else
		origin=0000;
		
end

/* �����֮�ǡ����׷��� */
always @(posedge clk_4Hz)	
begin

if(select)
begin

	/* ȫ���ܽ����� */
	if(state ==193)
		/* �Զ��ط� */
		state = 0;
	else
		/* ���ļ��� */
		state = state + 1'b1; 
	
	case(state)
		/* ��С�ڼ�� */
		/* 1 */
		0:											{high,med,low}='b000001100000;//��6
		1:					    					{high,med,low}='b000010000000;//��7
					
		/* 2 */
		2,3,4:									{high,med,low}='b000100000000;//��1
		5:											{high,med,low}='b000010000000;//��7
		6,7:                					{high,med,low}='b000100000000;//��1
		8,9:										{high,med,low}='b001100000000;//��3
					
		/* 3 */
		10,11,12,13,14,15:					{high,med,low}='b000010000000;//��7
		16,17:            					{high,med,low}='b000000110000;//��3
		
		/* 4 */		
		18,19,20:								{high,med,low}='b000001100000;//��6
		21:		 								{high,med,low}='b000001010000;//��5
		22,23:              	 				{high,med,low}='b000001100000;//��6
		24,25:									{high,med,low}='b000100000000;//��1
		
		/* 5 */
		26,27,28,29,30,31:					{high,med,low}='b000001010000;//��5   							
		32:				       				{high,med,low}='b000000100000;//��2
		33:			          				{high,med,low}='b000000110000;//��3
		
		/* 6 */
		34,35,36:				 				{high,med,low}='b000000111000;//��4
		37:					    				{high,med,low}='b000000110000;//��3
		38,39:					   			{high,med,low}='b000000111000;//��4
		40,41:				 					{high,med,low}='b000100000000;//��1
		
		/* 7 */
		42,43,44,45,46,47:      			{high,med,low}='b000000110000;//��3
		48,49:			    					{high,med,low}='b000100000000;//��1
		
		/* 8 */
		50,51,52:		       				{high,med,low}='b000010000000;//��7
		53,54,55:             				{high,med,low}='b000000111000;//��4
		56,57:									{high,med,low}='b000010000000;//��7
		
		/* 9 */
		58,59,60,61,62,63:					{high,med,low}='b000010000000;//��7
		64:					    				{high,med,low}='b000001100000;//��6
		65:				       				{high,med,low}='b000010000000;//��7
		
		/* 10 */
		66,67,68:	          				{high,med,low}='b000100000000;//��1
		69:					    				{high,med,low}='b000010000000;//��7
		70,71:			       				{high,med,low}='b000100000000;//��1
		72,73:			       				{high,med,low}='b001100000000;//��3
		
		/* 11 */
		74,75,76,77,78,79:					{high,med,low}='b000010000000;//��7
		80,81:			       				{high,med,low}='b000000110000;//��3
		
		/* 12 */
		82,83,84:    			 				{high,med,low}='b000001100000;//��6
		85:					    				{high,med,low}='b000000000101;//��5
		86,87:			       				{high,med,low}='b000001100000;//��6			
		88,89:                				{high,med,low}='b000100000000;//��1
		
		/* 13 */
		90,91,92,93,94,95:	 				{high,med,low}='b000001010000;//��5   							
		96:				       				{high,med,low}='b000000100000;//��2
		97:			          				{high,med,low}='b000000110000;//��3
		
		/* 14 */
		98,99:			 		 				{high,med,low}='b000000111000;//��4 
		100:					    				{high,med,low}='b000100000000;//��1
		101,102,103:							{high,med,low}='b000010000000;//��7
		104,105:					 				{high,med,low}='b000100000000;//��1
		
		/* 15 */
		106,107:					 				{high,med,low}='b001000000000;//��2
		108:						 				{high,med,low}='b001100000000;//��3
		109,110,111,112,113:					{high,med,low}='b000100000000;//��1
		
		/* 16 */
		114:										{high,med,low}='b000100000000;//��1
		115:		         			    	{high,med,low}='b000010000000;//��7			
		116:								 		{high,med,low}='b000001100000;//��6
		117:								 		{high,med,low}='b000001010000;//��5		
		118,119:								 	{high,med,low}='b000010000000;//��7
		120,121:								 	{high,med,low}='b000001010000;//��5
		
		/* 17 */
		122,123,124,125,126,127:			{high,med,low}='b000001100000;//��6
		128:					 					{high,med,low}='b000100000000;//��1
		129:						 				{high,med,low}='b001000000000;//��2
		
		/* 18 */
		130,131,132:    						{high,med,low}='b001100000000;//��3
		133:										{high,med,low}='b001000000000;//��2
		134,135:									{high,med,low}='b001100000000;//��3			
		136,137:            					{high,med,low}='b010000000000;//��5
		
		/* 19 */
		138,139,140,141,142,143:			{high,med,low}='b001000000000;//��2
		144,145:									{high,med,low}='b000001010000;//��5
		
		/* 20 */
		146,147,148:    						{high,med,low}='b000100000000;//��1
		149:										{high,med,low}='b000010000000;//��7
		150,151:									{high,med,low}='b000100000000;//��1
		152,153:									{high,med,low}='b001100000000;//��3
		
		/* 21 */
		154,155,156,157,158,159,160,161:	{high,med,low}='b000010000000;//��7
		
		/* 22 */
		162:										{high,med,low}='b000001100000;//��6
		163:										{high,med,low}='b000010000000;//��7
		164,165:									{high,med,low}='b000100000000;//��1
		166:										{high,med,low}='b000010000000;//��7
		167:										{high,med,low}='b000100000000;//��1
		168,169:									{high,med,low}='b001000000000;//��2
		
		/* 23 */
		170,171,172:							{high,med,low}='b000100000000;//��1	
		173,174,175,176,177:					{high,med,low}='b000001010000;//��5
		
		/* 24 */
		178,179:									{high,med,low}='b001010000000;//��4
		180,181:									{high,med,low}='b001100000000;//��3								
		182,183:									{high,med,low}='b001000000000;//��2
		184,185:									{high,med,low}='b000100000000;//��1
		
		/* 25 */
		186,187,188,189,190,191,192,193:	{high,med,low}='b001100000000;//��3	
	
	endcase

end

end

endmodule









